package my_pkg;
    import uvm_pkg::*;
    
    `include "uvm_macros.svh"
    `include "My_sequence_item.svh"
    `include "My_sequence.svh"
    `include "My_sequencer.svh"
    `include "My_driver.svh"
    `include "My_monitor.svh"
    `include "My_agent.svh"
    `include "My_subscriber.svh"
    `include "My_scoreboard.svh"
    `include "My_env.svh"
    `include "My_test.svh"
endpackage
